`include "CPU.v"

module tb;
    reg CLK, RESET;
    //output [31:0] PC;
    reg [31:0] INSTRUCTION ;
    //00000101_00000000_00000100_00000000 
   // 00001001_00000000_00000010_00000000               
   // 00000010_00000100_00000110_00000010
    wire WRITEENABLE;
    wire [2:0] ALUOP;
    wire COMPLEMENT_FLAG;
    wire IMMEDIATE_FALG;
	
    control_unit myctrlunit(INSTRUCTION,WRITEENABLE,ALUOP,COMPLEMENT_FLAG,IMMEDIATE_FALG);

    always begin
        CLK = 1; 
        $monitor($time,"INSTRUCTION=%b ,WRITEENABLE=%d ,ALUOP=%d ,COMPLEMENT_FLAG=%d,IMMEDIATE_FALG=%d",INSTRUCTION,WRITEENABLE,ALUOP,COMPLEMENT_FLAG,IMMEDIATE_FALG);
        #4 CLK = ~ CLK;
    end

    initial begin
        RESET =1;#4 RESET =0;
        #8 
        INSTRUCTION = 32'B00000101_00000000_00000100_00000000;//loadi 4 0x05
        #16
        INSTRUCTION = 32'B00001001_00000000_00000010_00000000;
       // $monitor($time,"INSTRUCTION=%b ,WRITEENABLE=%d ,ALUOP=%d ,COMPLEMENT_FLAG=%d,IMMEDIATE_FALG=%d\n",INSTRUCTION,WRITEENABLE,ALUOP,COMPLEMENT_FLAG,IMMEDIATE_FALG);
        #200 $finish;
    end

endmodule
