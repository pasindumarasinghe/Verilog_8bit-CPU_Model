
module cpu(PC, INSTRUCTION, CLK, RESET)
    
endmodule

module control_unit()

endmodule